--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package divisionPkg is

type divisionState is (Intial_state, Shift_state, Calculation_state, RemainderUPD_state, STOP);


end divisionPkg;

package body divisionPkg is

 
end divisionPkg;
